module debug_datos(
    input datos_adc,
    input datos_dac,
    input clock,
    output LED
    );


endmodule
